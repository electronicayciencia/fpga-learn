`timescale 1 ns/1 ns  // time-unit = 1 ns, precision = 10 ps

/*
 Now with a FSM. Send null-terminated string.

 Main top-level module

    PIN
    35  clock 24Mhz
    14  btn_b
    15  btn_a

 Logic ann. config for debug:
    45  Ch0  debug[0]
    11  Ch1  debug[1]
    44  Ch2  debug[2]
    43  Ch4  debug[3]
    10  Ch5  debug[4]
    42  Ch6  debug[5]
    46  Ch7  debug[6]
*/
module main_tb (
    input btn_a,
    input btn_b,
    input clk_i,
    output [6:0] debug
);


reg sys_clk = 0;

initial begin
	forever #333 sys_clk = ~sys_clk;
end


/*
    wire sys_clk; // slow clock for logic ann
    clkdiv Clkdiv1(
        .clk_i(clk_i),
        .clk_o(sys_clk)
    );
*/

    wire busy;
    wire start;
    wire restart;
    wire [3:0] address;
    wire [7:0] byte;

    /* Automatic restart */
    timer Timer1 (
        .clk_i(sys_clk),
        .clk_o(restart)
    );

    memory Mem(
        .clk_i(sys_clk),
        .addr_i(address),
        .data_o(byte)
    );

    baudclock UARTClk(
        .clk_i(sys_clk),
        .clk_o(uart_clk)
    );

    simpleUARTtx UART1 (
        .data(byte),
        .start(start),
        .clk(uart_clk),
        .busy(busy),
        .line(serial)
    );

    fsm FSM1 (
        .clk_i(sys_clk),
        .restart_i(restart),
        .byte_i(byte),
        .busy_i(busy),
        .start_o(start),
        .address_o(address)
    );
    




    assign debug[0] = restart;
    assign debug[1] = start;
    assign debug[2] = uart_clk;
    assign debug[3] = 0;
    assign debug[4] = serial;
    assign debug[5] = busy;
    assign debug[6] = sys_clk;

endmodule
module and_gate (
    input a, b,
    output o
);

assign o = a & b;

endmodule

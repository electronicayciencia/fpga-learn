module led (input btn, output led);

    assign led = btn;

endmodule


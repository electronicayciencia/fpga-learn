//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1N-LV1QN48C6/I5
//Device: GW1N-1
//Created Time: Sun Nov 07 14:14:47 2021

module chr_rom (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [9:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,ad[9:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_08 = 256'h006C6CFE6CFE6C6C0000000000006C6C00180018183C3C180000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000000C060600076CCDC76386C3800C6663018CCC6000030F80C78C07C30;
defparam prom_inst_0.INIT_RAM_0A = 256'h00003030FC3030000000663CFF3C660000603018181830600018306060603018;
defparam prom_inst_0.INIT_RAM_0B = 256'h0080C06030180C06003030000000000000000000FC0000006030300000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h0078CC0C380CCC7800FCCC60380CCC7800FC303030307030007CE6F6DECEC67C;
defparam prom_inst_0.INIT_RAM_0D = 256'h00303030180CCCFC0078CCCCF8C060380078CC0C0CF8C0FC001E0CFECC6C3C1C;
defparam prom_inst_0.INIT_RAM_0E = 256'h603030000030300000303000003030000070180C7CCCCC780078CCCC78CCCC78;
defparam prom_inst_0.INIT_RAM_0F = 256'h00300030180CCC78006030180C1830600000FC0000FC000000183060C0603018;
defparam prom_inst_0.INIT_RAM_10 = 256'h003C66C0C0C0663C00FC66667C6666FC00CCCCFCCCCC78300078C0DEDEDEC67C;
defparam prom_inst_0.INIT_RAM_11 = 256'h003E66CEC0C0663C00F06068786862FE00FE6268786862FE00F86C6666666CF8;
defparam prom_inst_0.INIT_RAM_12 = 256'h00E6666C786C66E60078CCCC0C0C0C1E007830303030307800CCCCCCFCCCCCCC;
defparam prom_inst_0.INIT_RAM_13 = 256'h00386CC6C6C66C3800C6C6CEDEF6E6C600C6C6D6FEFEEEC600FE6662606060F0;
defparam prom_inst_0.INIT_RAM_14 = 256'h0078CC1C70E0CC7800E6666C7C6666FC001C78DCCCCCCC7800F060607C6666FC;
defparam prom_inst_0.INIT_RAM_15 = 256'h00C6EEFED6C6C6C6003078CCCCCCCCCC00FCCCCCCCCCCCCC007830303030B4FC;
defparam prom_inst_0.INIT_RAM_16 = 256'h007860606060607800FE6632188CC6FE0078303078CCCCCC00C66C38386CC6C6;
defparam prom_inst_0.INIT_RAM_17 = 256'hFF0000000000000000000000C66C381000781818181818780002060C183060C0;
defparam prom_inst_0.INIT_RAM_18 = 256'h0078CCC0CC78000000DC66667C6060E00076CC7C0C7800000000000000183030;
defparam prom_inst_0.INIT_RAM_19 = 256'hF80C7CCCCC76000000F06060F0606C380078C0FCCC7800000076CCCC7C0C0C1C;
defparam prom_inst_0.INIT_RAM_1A = 256'h00E66C786C6660E078CCCC0C0C0C000C007830303070003000E66666766C60E0;
defparam prom_inst_0.INIT_RAM_1B = 256'h0078CCCCCC78000000CCCCCCCCF8000000C6D6FEFECC00000078303030303070;
defparam prom_inst_0.INIT_RAM_1C = 256'h00F80C78C07C000000F0606676DC00001E0C7CCCCC760000F0607C6666DC0000;
defparam prom_inst_0.INIT_RAM_1D = 256'h006CFEFED6C60000003078CCCCCC00000076CCCCCCCC000000183430307C3010;
defparam prom_inst_0.INIT_RAM_1E = 256'h001C3030E030301C00FC643098FC0000F80C7CCCCCCC000000C66C386CC60000;
defparam prom_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000DC7600E030301C3030E00018181800181818;

endmodule //chr_rom

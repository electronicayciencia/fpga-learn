module led (input i_btn, output o_led);

    assign o_led = i_btn;

endmodule


//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1N-LV1QN48C6/I5
//Device: GW1N-1
//Created Time: Tue Nov 09 14:02:13 2021

module text_ram (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [15:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [9:0] ada;
input [15:0] din;
input [9:0] adb;

wire [15:0] sdpb_inst_0_dout_w;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[15:0],dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 16;
defparam sdpb_inst_0.BIT_WIDTH_1 = 16;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E016170060706;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_02 = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_10 = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_12 = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_14 = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_1D = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_20 = 256'h072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_21 = 256'h072D072D072E072E072E072E072E072E072E072E072E072E072E072E072E072E;
defparam sdpb_inst_0.INIT_RAM_22 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_23 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_24 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_25 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_26 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_27 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_28 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_29 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_2A = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_2B = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_2C = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_2D = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_2E = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_2F = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_30 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_31 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_32 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_33 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_34 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_35 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_36 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_37 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_38 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_39 = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_3A = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_3B = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_3C = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_3D = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_3E = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;
defparam sdpb_inst_0.INIT_RAM_3F = 256'h072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D072D;

endmodule //text_ram

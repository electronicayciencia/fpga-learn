module and_gate (
    input i,
    output o
);

assign o = i;

endmodule
